`timescale 1ns/1ns
module osc_spice(
	dvddgo1,
	dvss ,
	id_en,
  od_clk 
);

   input dvddgo1, dvss, id_en;
   output od_clk;
   
endmodule // osc_spice
