* SPICE export by:  S-Edit 15.10
* Export time:      Fri Dec 16 10:44:13 2011
* Design:           rtest
* Cell:             carac_mos
* Interface:        schematic
* View:             schematic
* View type:        connectivity
* Export as:        top-level cell
* Export mode:      hierarchical
* Exclude empty cells: yes
* Exclude .model:   yes
* Exclude .end:     yes
* Exclude simulator commands:     yes
* Expand paths:     yes
* Wrap lines:       80 characters
* Root path:        \\VBOXSVR\aferret\virtualbox\tanner\sedit\rtest
* Exclude global pins:   yes
* Exclude instance locations: yes
* Control property name: SPICE

***** Top Level *****
CCLOAD ac_VD SUB cload
IID_AC VDD ac_VD DC id AC 0 0
VVALIM VDD SUB DC valim AC 0 0
VVDS_DC dc_VD dc_VS DC vds AC 0 0
VVG_AC ac_VG SUB DC vg AC 1 0
VVG_DC dc_VG SUB DC vg AC 0 0
VVS_AC ac_VS SUB DC vs AC 0 0
VVS_DC dc_VS SUB DC vs AC 0 0
XMN_AC ac_VD ac_VG ac_VS  SUB nmodel l=lngo1 w=wngo1 m=mngo1 nf=nfngo1 as='2*(wngo1/nfngo1*75e-9)+(nfngo1/2-1)*(wngo1/nfngo1*100e-9)' 
+ad='0.5*wngo1*100n' ps='2*(2*(wngo1/nfngo1+75e-9)+(nfngo1/2-1)*(wngo1/nfngo1+100e-9))' 
+pd='2*(0.5*wngo1+100n)' sa='(1/nfngo1)*(nfngo1*75e-9+0.5*(nfngo1*(nfngo1-1))*(lngo1+100e-9))' 
+sb='(1/nfngo1)*(nfngo1*75e-9+0.5*(nfngo1*(nfngo1-1))*(lngo1+100e-9))'
XMN_DC dc_VD dc_VG dc_VS  SUB nmodel l=ln w='wnf*nnf' m=mn nf=nnf


