
  --Write register
  isolation_n           <= control_reg_o(0);
  TxClkPolarity         <= control_reg_o(1);
  TxPisoSelTxSync       <= control_reg_o(2);
  TxCtrlMain            <= control_reg_o(6 downto 3);
  TxCtrlPre             <= control_reg_o(10 downto 7);
  TxCtrlTest            <= control_reg_o(14 downto 11);
  TxDataSelect          <= control_reg_o(15);
  TxDciPup              <= control_reg_o(16);
  TxPisoDivInit         <= control_reg_o(20 downto 17);
  TxPisoReset           <= control_reg_o(21);
  TxPisoSelDiv          <= control_reg_o(22);
  TxPreEmph             <= control_reg_o(23);
  TxPup                 <= control_reg_o(24);
  TxRtrim               <= control_reg_o(29 downto 25);
  TxRxLpbkSelect        <= control_reg_o(30);
  TxTestLpbk            <= control_reg_o(31);
  TxTestPcsEn           <= control_reg_o(32);
  cmn_bias_on           <= control_reg_o(33);
  cmn_dci_dc            <= control_reg_o(35 downto 34);
  cmn_dci_prog          <= control_reg_o(40 downto 36);
  sx_vco_cc             <= control_reg_o(42 downto 41);
  sx_PupDco_Out         <= control_reg_o(43);
  TxClkSync_inv         <= control_reg_o(44);
  cmn_spare             <= control_reg_o(63 downto 48);
  -- 2nd reg
  sx_DivN               <= control_reg_o(69 downto 64);
  sx_DpllAlpha          <= control_reg_o(72 downto 70);
  sx_DpllBeta           <= control_reg_o(75 downto 73);
  sx_DpllOpenLoop       <= control_reg_o(84 downto 76);
  sx_DpllReset          <= control_reg_o(85);
  sx_Dpll_Fcw           <= control_reg_o(91 downto 86);
  sx_Dpll_FiltMux       <= control_reg_o(92);
  sx_Dpll_VarDem        <= control_reg_o(93);
  sx_FrefDciGnd         <= control_reg_o(94);
  sx_FrefDciProg50      <= control_reg_o(99 downto 95);
  sx_FrefDciVdd         <= control_reg_o(100);
  sx_FrefPup            <= control_reg_o(101);
  sx_LoExtDciGnd        <= control_reg_o(102);
  sx_LoExtDciProg50     <= control_reg_o(107 downto 103);
  sx_LoExtDciVdd        <= control_reg_o(108);
  sx_LoExtPup           <= control_reg_o(109);
  sx_LoSrcMux           <= control_reg_o(110);
  sx_PupLoRx            <= control_reg_o(111);
  sx_PupLoTx            <= control_reg_o(112);
  sx_PupRefOut          <= control_reg_o(113);
  sx_RxDiv              <= control_reg_o(116 downto 114);
--  sx_TxDiv              <= control_reg_o(119 downto 117); " chevauchement de 2 registres "
  sx_TxDiv              <= control_reg_o(274 downto 272);
  sx_filter_size        <= control_reg_o(126 downto 118);
  sx_pll_typ            <= control_reg_o(127);
  -- 3rd and 4th regs
  rx_bias_off           <= control_reg_o(130 downto 128);
  rx_cdr_en             <= control_reg_o(131);
  rx_cdr_filt_openloop  <= control_reg_o(144 downto 132);
  rx_cdr_filta          <= control_reg_o(147 downto 145);
  -- 148 missing
  rx_cdr_filtb          <= control_reg_o(151 downto 149);
  rx_cdr_filtc          <= control_reg_o(154 downto 152);
  rx_cdr_rst            <= control_reg_o(155);
  rx_cdr_sel_openloop   <= control_reg_o(156);
  rx_cdr_var_dem        <= control_reg_o(157);
  rx_clk_dela           <= control_reg_o(165 downto 158);
  rx_clk_delb           <= control_reg_o(173 downto 166);
  rx_clk_en             <= control_reg_o(174);
  rx_clk_sel            <= control_reg_o(175);
  -- 176 missing
  rx_cmp_aux_en         <= control_reg_o(177);
  rx_cmp_off            <= control_reg_o(178);
  rx_cmp_thhigh         <= control_reg_o(183 downto 179);
  rx_cmp_thlow          <= control_reg_o(188 downto 184);
  rx_dfe_coef1          <= control_reg_o(193 downto 189);
  rx_dfe_coef2          <= control_reg_o(198 downto 194);
  rx_dfe_en             <= control_reg_o(199);
  rx_ff_gain1           <= control_reg_o(201 downto 200);
  rx_ff_gain2           <= control_reg_o(203 downto 202);
  rx_ff_off             <= control_reg_o(206 downto 204);
  rx_ff_setresc         <= control_reg_o(209 downto 207);
  rx_ff_setresr         <= control_reg_o(212 downto 210);
  rx_in_dccouple        <= control_reg_o(213);
  rx_in_load50          <= control_reg_o(218 downto 214);
  rx_in_load100k        <= control_reg_o(220 downto 219);
  rx_in_ref50           <= control_reg_o(222 downto 221);
--  rx_loopback1_en       <= control_reg_o(223);
  rx_loopback2_rx2tx_en <= control_reg_o(224);
  rx_loopback2_tx2rx_en <= control_reg_o(225);
-- rxout0 <= control_reg_o(226);
-- rxout1 <= control_reg_o(227);
  rx_sel_data           <= control_reg_o(228);
  rx_sel_test           <= control_reg_o(233 downto 229);
  rx_sipo_aux_sel       <= control_reg_o(235 downto 234);
  rx_sipo_en            <= control_reg_o(236);
  rx_sipo_invdata       <= control_reg_o(237);
  rx_sipo_n             <= control_reg_o(241 downto 238);
  rx_sipo_rst           <= control_reg_o(242);
  rx_vref_bypass        <= control_reg_o(243);
  rx_sipo_seldiv        <= control_reg_o(244);
  rx_cdr_sel_data       <= control_reg_o(247 downto 245);
  rx_cdr_sel_clk        <= control_reg_o(250 downto 248);
  -- 5th reg => spare bits and thermal sensor
  tx_spare              <= control_reg_o(271 downto 256);
  sx_spare              <= control_reg_o(287 downto 272);
  rx_spare              <= control_reg_o(303 downto 288);
  th_enad               <= control_reg_o(304);
  th_envref             <= control_reg_o(305);
  th_enbgr              <= control_reg_o(306);
  th_stn                <= control_reg_o(307);
  th_tmod               <= control_reg_o(308);
  th_itcl               <= control_reg_o(310 downto 309);
  th_spare              <= control_reg_o(318 downto 311);
  -- 6th and 7th regs => PRBS control

  --status_i((2*64)+19 downto (2*64)+9) <= th_dataready & th_data;
  --status_i((6*64)-1 downto (2*64)+20) <= (others => '0');
  --rx_err_cnt_o      => status_i((1*64)-1 downto 0*64),
  --rx_cnt_o          => status_i((2*64)-1 downto 1*64),
  --prbs_config_sta_o => status_i((7*64)-1 downto 6*64),
  --prbs_config_ctl_i => control_reg_o((6*64)-1 downto 5*64)
  -- Modified affectation & number
  -- In order to ease script, different status for Hash Table & read ...
  -- Read Register
  status_i(147 downto 137) <= th_dataready & th_data;
  status_i(383 downto 148) <= null ;
  status_i(63 downto 0) <= rx_err_cnt_o;
  status_i(127 downto 64) <= rx_cnt_o;
  status_i(447 downto 384) <= prbs_config_sta_o;
  control_reg_o(383 downto 320) <= prbs_config_ctl_i; 
  regtest(383) <= prbs_config_test_i; 

  control_rst_val(218 downto 214) <= "10000";  -- rx_in_load50          
  control_rst_val(222 downto 221) <= "10";  -- rx_in_ref50           
  control_rst_val(213)            <= '1';  -- rx_in_dccouple        
  control_rst_val(220 downto 219) <= "11";  -- rx_in_load100k        
  control_rst_val(201 downto 200) <= "10";  -- rx_ff_gain1           
  control_rst_val(203 downto 202) <= "01";  -- rx_ff_gain2           
  control_rst_val(209 downto 207) <= "011";  -- rx_ff_setresc         
  control_rst_val(212 downto 210) <= "011";  -- rx_ff_setresr         
  control_rst_val(174)            <= '1';  -- rx_clk_en             
  control_rst_val(241 downto 238) <= "1000";  -- rx_sipo_n             
  control_rst_val(244)            <= '1';  -- rx_sipo_seldiv        
  control_rst_val(144 downto 132) <= "0010111011100";  -- rx_cdr_filt_openloop  
  control_rst_val(147 downto 145) <= "010";  -- rx_cdr_filta          
  control_rst_val(151 downto 149) <= "011";  -- rx_cdr_filtb          
  control_rst_val(154 downto 152) <= "010";  -- rx_cdr_filtc          
  control_rst_val(112)            <= '1';  -- sx_PupLoTx            
  control_rst_val(110)            <= '1';  -- sx_LoSrcMux           
  control_rst_val(111)            <= '1';  -- sx_PupLoRx            
  control_rst_val(75 downto 73)   <= "010";  -- sx_DpllBeta           
  control_rst_val(126 downto 118) <= "111111111";  -- sx_filter_size        
  control_rst_val(91 downto 86)   <= "011001";  -- sx_Dpll_Fcw           
  control_rst_val(69 downto 64)   <= "000111";  -- sx_DivN               
  control_rst_val(107 downto 103) <= "10000";  -- sx_LoExtDciProg50     
  control_rst_val(108)            <= '1';  -- sx_LoExtDciVdd        
  control_rst_val(99 downto 95)   <= "10000";  -- sx_FrefDciProg50      
  control_rst_val(101)            <= '1';  -- sx_FrefPup            
  control_rst_val(100)            <= '1';  -- sx_FrefDciVdd         
  control_rst_val(127)            <= '1';  -- sx_pll_typ            
-- mike modif: control_rst_val(20 downto 17) 1111 => 1000  "erreur dans le fichier xls"
  control_rst_val(20 downto 17)   <= "1000";  -- TxPisoDivInit         
  control_rst_val(24)             <= '1';  -- TxPup                 
  control_rst_val(6 downto 3)     <= "1000";  -- TxCtrlMain            
  control_rst_val(10 downto 7)    <= "0001";  -- TxCtrlPre             
  control_rst_val(16)             <= '1';  -- TxDciPup              
  control_rst_val(29 downto 25)   <= "01111";  -- TxRtrim               
  control_rst_val(33)             <= '1';  -- cmn_bias_on           
  control_rst_val(35 downto 34)   <= "10";  -- cmn_dci_dc            
  control_rst_val(40 downto 36)   <= "10000";  -- cmn_dci_prog          
-- mike modif: ontrol_rst_val(42 downto 41) 00 => 01
  control_rst_val(42 downto 41)   <= "01";  -- sx_vco_cc
  control_rst_val(305)            <= '1';  -- th_envref             
  control_rst_val(306)            <= '1';  -- th_enbgr              
  control_rst_val(318 downto 311) <= "00001010";  -- th_spare

